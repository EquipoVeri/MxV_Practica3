module FSM_MxV_Control(
);

endmodule
